library verilog;
use verilog.vl_types.all;
entity UC_PLUS_TIMER_vlg_sample_tst is
    port(
        ADD             : in     vl_logic;
        \AND\           : in     vl_logic;
        clk             : in     vl_logic;
        flagN           : in     vl_logic;
        flagZ           : in     vl_logic;
        HLT             : in     vl_logic;
        JMP             : in     vl_logic;
        JN              : in     vl_logic;
        JZ              : in     vl_logic;
        LDA             : in     vl_logic;
        NOP             : in     vl_logic;
        \NOT\           : in     vl_logic;
        \OR\            : in     vl_logic;
        Reset           : in     vl_logic;
        STA             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end UC_PLUS_TIMER_vlg_sample_tst;
