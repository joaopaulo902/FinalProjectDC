library verilog;
use verilog.vl_types.all;
entity AC_vlg_vec_tst is
end AC_vlg_vec_tst;
