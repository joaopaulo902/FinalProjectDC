library verilog;
use verilog.vl_types.all;
entity UC_PLUS_TIMER_vlg_vec_tst is
end UC_PLUS_TIMER_vlg_vec_tst;
