library verilog;
use verilog.vl_types.all;
entity flagLogic_vlg_vec_tst is
end flagLogic_vlg_vec_tst;
