library verilog;
use verilog.vl_types.all;
entity Mux8bit_vlg_vec_tst is
end Mux8bit_vlg_vec_tst;
