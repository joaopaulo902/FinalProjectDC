library verilog;
use verilog.vl_types.all;
entity NEANDER_vlg_vec_tst is
end NEANDER_vlg_vec_tst;
