library verilog;
use verilog.vl_types.all;
entity feqDiv_vlg_vec_tst is
end feqDiv_vlg_vec_tst;
